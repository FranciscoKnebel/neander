--
-- Authors: Francisco Paiva Knebel
--				Gabriel Alexandre Zillmer
--
-- Universidade Federal do Rio Grande do Sul
-- Instituto de Inform�tica
-- Sistemas Digitais
-- Prof. Fernanda Lima Kastensmidt
--
-- Create Date:    09:49:46 05/03/2016 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity neander is
end neander;

architecture Behavioral of neander is
begin

	

end Behavioral;

